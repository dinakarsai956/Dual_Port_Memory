`include "dual_port_memory_latency.sv"
`include "hamming_encoder.sv"
`include "hamming_decoder.sv"
`include "multi_bank_memory.sv"
