//`include"packet.sv"
`include"transaction.sv"
`include"interface.sv"
`include"generator.sv"
`include"driver.sv"
`include"monitor.sv"
`include"reference.sv"
`include"scoreboard.sv"
`include"environment.sv"

